//Block Code
parameter ACORTEX_BLK               = 4'd0;
parameter VCORTEX_BLK               = 4'd1;
parameter FGYRUS_BLK                = 4'd2;
