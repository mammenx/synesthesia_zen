//Block Code
parameter VCORTEX_GPU_CODE      =    4'd0;
parameter VCORTEX_VGA_CODE      =    4'd1;

//Grapheme register addresses
parameter VCORTEX_GPU_CONTROL_REG_ADDR      = 8'd0;
parameter VCORTEX_GPU_STATUS_REG_ADDR       = 8'd1;
parameter VCORTEX_GPU_JOB_BFFR_0_REG_ADDR   = 8'd2;
parameter VCORTEX_GPU_JOB_BFFR_1_REG_ADDR   = 8'd3;
parameter VCORTEX_GPU_JOB_BFFR_2_REG_ADDR   = 8'd4;
parameter VCORTEX_GPU_JOB_BFFR_3_REG_ADDR   = 8'd5;
parameter VCORTEX_GPU_JOB_BFFR_4_REG_ADDR   = 8'd6;
parameter VCORTEX_GPU_JOB_BFFR_5_REG_ADDR   = 8'd7;
parameter VCORTEX_GPU_JOB_BFFR_6_REG_ADDR   = 8'd8;
parameter VCORTEX_GPU_JOB_BFFR_7_REG_ADDR   = 8'd9;
